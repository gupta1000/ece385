module testbench();

timeunit 10ns;	// Half clock cycle at 50 MHz
			// This is the amount of time represented by #1
timeprecision 1ns;

// These signals are internal because the processor will be
// instantiated as a submodule in testbench.
logic Clk = 0;
logic Reset, Run, Continue, CE, UB, LB, OE, WE;
logic [15:0] S, IR;
logic [11:0] LED;
logic [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, HEX6, HEX7;
logic [19:0] ADDR;
wire [15:0] Data;

// Instantiating the DUT
// Make sure the module and signal names match with those in your design
lab6_toplevel lab6(.*);

// Toggle the clock
// #1 means wait for a delay of 1 timeunit
always begin : CLOCK_GENERATION
#1 Clk = ~Clk;
end

initial begin: CLOCK_INITIALIZATION
    Clk = 0;
end

// Testing begins here
// The initial block is not synthesizable
// Everything happens sequentially inside an initial block
// as in a software program
initial begin: TEST_VECTORS

	// init the state of the essential signals in simulation
	Reset = 0;
	Run = 1;
	Continue = 1;

	// set switches to a program (bubblesort)
	S = 16'h005a;

	#2 Reset = 1;

	// start program
	#2 Run = 0;
	#2 Run = 1;

	#20 Continue = 0;

	// repeatedly press and release continue
	for(int i = 0; i < 10; i++)
	begin
		#2 Continue = 0;
		#2 Continue = 1;
	end

	// set switches to another value (sort)
	#2 S = 16'h0002;

	// repeatedly press continue
	for(int i = 0; i < 40000; i++)
	begin
		#2 Continue = 0;
		#2 Continue = 1;
	end

	// set switches to another value (display values)
	#2 S = 16'h0003;

	// repeatedly press continue
	for(int i = 0; i < 40000; i++)
	begin
		#2 Continue = 0;
		#2 Continue = 1;
	end

end
endmodule
